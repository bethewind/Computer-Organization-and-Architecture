module notgate(
    input x,
    output p
);

assign p = ~x;
endmodule

